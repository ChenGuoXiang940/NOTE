library verilog;
use verilog.vl_types.all;
entity ENCODER4_2_vlg_vec_tst is
end ENCODER4_2_vlg_vec_tst;
