library verilog;
use verilog.vl_types.all;
entity RELATIONAL_vlg_vec_tst is
end RELATIONAL_vlg_vec_tst;
