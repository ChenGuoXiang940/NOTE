library verilog;
use verilog.vl_types.all;
entity test is
    port(
        I               : in     vl_logic_vector(8 downto 0);
        pe              : out    vl_logic
    );
end test;
