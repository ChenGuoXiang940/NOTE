library verilog;
use verilog.vl_types.all;
entity MUL2_1 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        S               : in     vl_logic;
        F               : out    vl_logic
    );
end MUL2_1;
