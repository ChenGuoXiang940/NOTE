library verilog;
use verilog.vl_types.all;
entity DUPLICATION_vlg_vec_tst is
end DUPLICATION_vlg_vec_tst;
