library verilog;
use verilog.vl_types.all;
entity AND_GATE_vlg_vec_tst is
end AND_GATE_vlg_vec_tst;
