library verilog;
use verilog.vl_types.all;
entity PRIORITY_vlg_vec_tst is
end PRIORITY_vlg_vec_tst;
