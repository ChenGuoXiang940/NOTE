library verilog;
use verilog.vl_types.all;
entity BITWISE_vlg_vec_tst is
end BITWISE_vlg_vec_tst;
