library verilog;
use verilog.vl_types.all;
entity MUL3_1_vlg_vec_tst is
end MUL3_1_vlg_vec_tst;
