library verilog;
use verilog.vl_types.all;
entity DECODER3_5_vlg_vec_tst is
end DECODER3_5_vlg_vec_tst;
