library verilog;
use verilog.vl_types.all;
entity MUL2_1_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MUL2_1_vlg_check_tst;
