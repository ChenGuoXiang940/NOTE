library verilog;
use verilog.vl_types.all;
entity D_FF2_vlg_vec_tst is
end D_FF2_vlg_vec_tst;
