library verilog;
use verilog.vl_types.all;
entity ENCODER4_2_vlg_check_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ENCODER4_2_vlg_check_tst;
