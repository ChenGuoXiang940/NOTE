library verilog;
use verilog.vl_types.all;
entity DEMUL1_4_vlg_vec_tst is
end DEMUL1_4_vlg_vec_tst;
