library verilog;
use verilog.vl_types.all;
entity LOGICAL_vlg_vec_tst is
end LOGICAL_vlg_vec_tst;
