library verilog;
use verilog.vl_types.all;
entity CONCATENATION_vlg_vec_tst is
end CONCATENATION_vlg_vec_tst;
