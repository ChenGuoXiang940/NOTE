library verilog;
use verilog.vl_types.all;
entity DECODER3_8_vlg_vec_tst is
end DECODER3_8_vlg_vec_tst;
