library verilog;
use verilog.vl_types.all;
entity MUL2_1_vlg_vec_tst is
end MUL2_1_vlg_vec_tst;
